library verilog;
use verilog.vl_types.all;
entity tb_float_conv_sv_unit is
end tb_float_conv_sv_unit;
