`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mf2iq8JtkesW284ST3Pyb2vw5SJXbSFCf+xCpU2+/pSBqtPkej1Bbqdi0TuU7IEo
uetIn8AuRD2twaCOiJq9gA2zashA9bferq28VllI2RAqAx30WzHeZmpDRLEW1gJG
EKcNIunLuQ3KOQ+TYrFP1w==
`protect END_PROTECTED
